----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/23/2025 05:55:26 PM
-- Design Name: 
-- Module Name: eth_top - rtl
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
-- eth_top.vhd will contain:
--      - eth_wishbone (?) (may replace with some kind of PCIe interface)
--      - eth_registers.vhd
--      - eth_rxethmac.vhd
--      - eth_macstatus.vhd
--      - eth_txethmac.vhd
--      - eth_maccontrol.vhd
--      - eth_miim.vhd
----------------------------------------------------------------------------------


library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity eth_top is
--  Port ( );
end eth_top;

architecture rtl of eth_top is

begin


end rtl;
